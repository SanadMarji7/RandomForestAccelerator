library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use std.textio.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;

entity DT_memory is
  Port (
        tree_num : in integer;
        currentNode : in std_logic_vector;
        allinf : out std_logic_vector(19 downto 0)
        );
end DT_memory;

architecture Behavioral of DT_memory is
--2-dimensional array used to store all information needed for all the decision trees in the random forest.
-- function InitRamFromFile below is used to read data stream from .data file generated by the python code(in Github)
--and store the data stream in the array. there are a total of 10 data chunks within the .data file
--each one of the 10 data chunks can hold 1-15 20-bit data streams each representing information of a node.
    type mem is array(0 to 9, 0 to 14) of std_logic_vector(19 downto 0);
   
    impure function InitRamFromFile (RamFileName : in string) return mem is
    file RamFile : text is in RamFileName;
    variable RamFileLine : line;
    variable RAM : mem;
    begin
        L1 : for i in 0 to 9 loop
            L2 : for j in 0 to 14 loop
                readline(RamFile, RamFileLine);
                if RamFileLine'length < 4 then
                    exit L2;
                else
                    read(RamFileLine, RAM(i,j));       
                end if;
            end loop;
        end loop;
        return RAM;   
   end function;
   
   --function InitRamFromFile called and the return value stored in signal RAM
   signal RAM : mem := InitRamFromFile("/home/marji/Desktop/Fachprojekt/DT_Data/randomForest.data");
begin
    -- data stream of each node is fetched.
    allinf <= RAM(tree_num, to_integer(unsigned(currentNode)));

end Behavioral;
