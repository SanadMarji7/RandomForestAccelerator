--10 instances of the DT component are called within the Random_Forest_accelerator design, each given a unique tree_number and the same sl, sw, pl, pw
--values to calculate their decisions simultaniously. this design shows how each decision is calculated in more detail.
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use std.textio.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;

--entity of design has:
--5 inputs: tree_number --> used for memory access, sl, sw, pl, pw --> used for calculating decision
--1 output: class_out --> contains final decision of decision tree.
entity DT is
    port(
    tree_number : in integer;
    sepal_length : in std_logic_vector(3 downto 0); 
    sepal_width : in std_logic_vector(3 downto 0); 
    petal_length : in std_logic_vector(3 downto 0); 
    petal_width : in std_logic_vector(3 downto 0); 
    class_out : out std_logic_vector(3 downto 0) 
    
    );
end DT;

architecture Behavioral of DT is
--2-dimensional array used to store all information needed for all the decision trees in the random forest.
-- function InitRamFromFile below is used to read data stream from .data file generated by the python code(in Github)
--and store the data stream in the array. there are a total of 10 data chunks within the .data file
--each one of the 10 data chunks can hold 1-15 20-bit data streams each representing information of a node.
   type mem is array(0 to 9, 0 to 14) of std_logic_vector(19 downto 0);
   
    impure function InitRamFromFile (RamFileName : in string) return mem is
    file RamFile : text is in RamFileName;
    variable RamFileLine : line;
    variable RAM : mem;
    begin
        L1 : for i in 0 to 9 loop
            L2 : for j in 0 to 14 loop
                readline(RamFile, RamFileLine);
                if RamFileLine'length < 4 then
                    exit L2;
                else
                    read(RamFileLine, RAM(i,j));       
                end if;
            end loop;
        end loop;
        return RAM;   
   end function;
   
   --function InitRamFromFile called and the return value stored in signal RAM
   signal RAM : mem := InitRamFromFile("/home/marji/Desktop/Fachprojekt/DT_Data/randomForest.data");

        
--use of component node within the decision tree architecture
    component node is
    port(
        all_info : in std_logic_vector(19 downto 0);
        feature_to_compare : in std_logic_vector(3 downto 0);
        next_node : out std_logic_vector(3 downto 0);
        current_node : in std_logic_vector(3 downto 0)
    );
    end component;
    
    signal currentNode, nextNode1, nextNode2, nextNode3 : std_logic_vector(3 downto 0);
    signal f1, f2, f3 : std_logic_vector(3 downto 0);
    signal allinf0, allinf1, allinf2, allinf3 : std_logic_vector(19 downto 0);
     
     --the blelow getFeature function takes one input and returns the feature to be used within the comparator to calculate the decision.
     --whenever feature given within parameter is:
     --0000=>sepal length must be used as feature to compare
     --0001=>sepal width must be used as feature to compare
     --0010=>petal length must be used as feature to compare
     --0011=>petal width must be used as feature to compare
     impure function getFeature (a : std_logic_vector) return std_logic_vector is 
     begin
        if a = "0000" then
            return sepal_length;
        elsif a = "0001" then
            return sepal_width;
        elsif a = "0010" then
            return petal_length;
        elsif a = "0011" then
            return petal_width;
        else return "0000";
        end if;
     end getFeature;
     
     --getInfo fetches the information of one node (20 bit std_logic_vector) it uses tree_number to fetch correct address as well.
     impure function getInfo (z : std_logic_vector) return std_logic_vector is
     variable addr : integer;
     begin
        addr := to_integer(unsigned(z));
        return RAM(tree_number, addr);
     end getInfo;

begin
    --the design must always start with current node 0(root node) which has first address in data file
    --20 bit-data of each node is fetched using the getInfo function
    --3 instances of the component node are created since there is a max_depth of 3, each instance returns the next node(either left or right child)
    --at the end we read the class from the last node the design has reached
     currentNode <= "0000";
     allinf0 <= getInfo(currentNode);
     f1 <= getFeature(allinf0(15 downto 12));
     instance_node_1 : node port map(all_info => allinf0, feature_to_compare => f1, next_node => nextNode1, current_node => currentNode);
     
     
     allinf1 <= getInfo(nextNode1);
     f2 <= getFeature(allinf1(15 downto 12)) after 1ns;
     instance_node_2 : node port map(all_info => allinf1, feature_to_compare => f2, next_node => nextNode2, current_node => nextNode1);
     
     allinf2 <= getInfo(nextNode2);
     f3 <= getFeature(allinf2(15 downto 12)) after 2ns;
     instance_node_3 : node port map(all_info => allinf2, feature_to_compare => f3, next_node => nextNode3, current_node => nextNode2);
     
     class_out <= getInfo(nextNode3)(3 downto 0);
     
end Behavioral;
